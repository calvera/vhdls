package crystal_pkg is
	constant crystal_hz: positive := 50_000_000;
end package;
